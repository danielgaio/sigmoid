// --------------------------------------------------------------------------------------------
// Nome do modulo: sigmoid
// Entradas: x = valor real negativo ou positivo
// Saidas: y = valor real negativo ou positivo
// Descriçao: Implementaçao de funçao sigmoid no intervalo [-7, 7]
// --------------------------------------------------------------------------------------------


module sigmoid(x, y);
	input signed [15:0]x;
	output reg signed [15:0]y;
	
	
	always @ (x) begin
		case (x)
		
			16'b1001_000000000000 : y <= 16'b0000_000000000000;					// if x == -7 then y = 0
			16'b1010_100000000000 : y <= 16'b0000_000000000110;
			16'b1010_000000000000 : y <= 16'b0000_000000001010;
			16'b1011_100000000000 : y <= 16'b0000_000000010001;
			16'b1011_000000000000 : y <= 16'b0000_000000011011;
			16'b1100_100000000000 : y <= 16'b0000_000000101101;
			16'b1100_000000000000 : y <= 16'b0000_000001001010;
			16'b1101_100000000000 : y <= 16'b0000_000001111000;
			16'b1101_000000000000 : y <= 16'b0000_000011000010;
			16'b1110_100000000000 : y <= 16'b0000_000101000010;
			16'b1110_000000000000 : y <= 16'b0000_000111101000;
			16'b1111_100000000000 : y <= 16'b0000_001011101011;
			16'b1111_000000000000 : y <= 16'b0000_010001001110;
			16'b0000_100000000000 : y <= 16'b0000_011000001010;
			16'b0000_000000000000 : y <= 16'b0000_100000000000;
			16'b0000_100000000000 : y <= 16'b0000_100111110110;
			16'b0001_000000000000 : y <= 16'b0000_101110110010;
			16'b0001_100000000000 : y <= 16'b0000_110100010101;
			16'b0010_000000000000 : y <= 16'b0000_111000011000;
			16'b0010_100000000000 : y <= 16'b0000_111011001001;
			16'b0011_000000000000 : y <= 16'b0000_111100111110;
			16'b0011_100000000000 : y <= 16'b0000_111110001000;
			16'b0100_000000000000 : y <= 16'b0000_111110110110;
			16'b0100_100000000000 : y <= 16'b0000_111111010011;
			16'b0101_000000000000 : y <= 16'b0000_111111100101;
			16'b0101_100000000000 : y <= 16'b0000_111111101111;
			16'b0110_000000000000 : y <= 16'b0000_111111110110;
			16'b0110_100000000000 : y <= 16'b0000_111111111010;
			16'b0111_000000000000 : y <= 16'b0001_000000000000;					// if x == 7 then y = 1
			default : begin
				if (x[15] == 1) 	y <= 16'b0000_000000000000;
				else 					y <= 16'b0001_000000000000;
			end
			
		endcase
	end
		

endmodule
